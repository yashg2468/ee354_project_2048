module tile_rom_4
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==10'b0000000000)) color_data = 12'b110111011011;
		if(({row_reg, col_reg}==10'b0000000001)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0000000010)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0000000011)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}>=10'b0000000100) && ({row_reg, col_reg}<10'b0000000110)) color_data = 12'b111111110111;
		if(({row_reg, col_reg}>=10'b0000000110) && ({row_reg, col_reg}<10'b0000001100)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}>=10'b0000001100) && ({row_reg, col_reg}<10'b0000001111)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}>=10'b0000001111) && ({row_reg, col_reg}<10'b0000011001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0000011001)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}>=10'b0000011010) && ({row_reg, col_reg}<10'b0000011100)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0000011100)) color_data = 12'b111111100111;

		if(({row_reg, col_reg}==10'b0000011101)) color_data = 12'b110111000100;
		if(({row_reg, col_reg}==10'b0000100000)) color_data = 12'b111011101100;
		if(({row_reg, col_reg}==10'b0000100001)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0000100010)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}>=10'b0000100011) && ({row_reg, col_reg}<10'b0000100110)) color_data = 12'b111111110111;
		if(({row_reg, col_reg}>=10'b0000100110) && ({row_reg, col_reg}<10'b0000111100)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0000111100)) color_data = 12'b111011010110;

		if(({row_reg, col_reg}==10'b0000111101)) color_data = 12'b110011000100;
		if(({row_reg, col_reg}==10'b0001000000)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0001000001)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0001000010)) color_data = 12'b111011010111;
		if(({row_reg, col_reg}==10'b0001000011)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}>=10'b0001000100) && ({row_reg, col_reg}<10'b0001001000)) color_data = 12'b110011000101;
		if(({row_reg, col_reg}>=10'b0001001000) && ({row_reg, col_reg}<10'b0001001010)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}==10'b0001001010)) color_data = 12'b110111000100;
		if(({row_reg, col_reg}>=10'b0001001011) && ({row_reg, col_reg}<10'b0001010011)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}>=10'b0001010011) && ({row_reg, col_reg}<10'b0001010110)) color_data = 12'b110011000101;
		if(({row_reg, col_reg}>=10'b0001010110) && ({row_reg, col_reg}<10'b0001011001)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}>=10'b0001011001) && ({row_reg, col_reg}<10'b0001011011)) color_data = 12'b110011000101;
		if(({row_reg, col_reg}==10'b0001011011)) color_data = 12'b110011000100;
		if(({row_reg, col_reg}==10'b0001011100)) color_data = 12'b101010100011;

		if(({row_reg, col_reg}==10'b0001011101)) color_data = 12'b101010100010;
		if(({row_reg, col_reg}==10'b0001100000)) color_data = 12'b111011101000;
		if(({row_reg, col_reg}==10'b0001100001)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==10'b0001100010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b0001100011) && ({row_reg, col_reg}<10'b0001100101)) color_data = 12'b110111000110;
		if(({row_reg, col_reg}>=10'b0001100101) && ({row_reg, col_reg}<10'b0001101000)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0001101000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0001101001) && ({row_reg, col_reg}<10'b0001101011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0001101011) && ({row_reg, col_reg}<10'b0001101110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0001101110) && ({row_reg, col_reg}<10'b0001110000)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}>=10'b0001110000) && ({row_reg, col_reg}<10'b0001110011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0001110011) && ({row_reg, col_reg}<10'b0001110101)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0001110101) && ({row_reg, col_reg}<10'b0001111000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0001111000)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b0001111001) && ({row_reg, col_reg}<10'b0001111011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0001111011)) color_data = 12'b101111000100;

		if(({row_reg, col_reg}>=10'b0001111100) && ({row_reg, col_reg}<10'b0010000000)) color_data = 12'b100110100010;
		if(({row_reg, col_reg}==10'b0010000000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0010000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0010000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0010000011)) color_data = 12'b110111000110;
		if(({row_reg, col_reg}>=10'b0010000100) && ({row_reg, col_reg}<10'b0010000110)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}>=10'b0010000110) && ({row_reg, col_reg}<10'b0010001000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0010001000) && ({row_reg, col_reg}<10'b0010001100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0010001100) && ({row_reg, col_reg}<10'b0010001110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0010001110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0010001111)) color_data = 12'b111111000101;
		if(({row_reg, col_reg}>=10'b0010010000) && ({row_reg, col_reg}<10'b0010010011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0010010011) && ({row_reg, col_reg}<10'b0010010101)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0010010101) && ({row_reg, col_reg}<10'b0010011000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0010011000) && ({row_reg, col_reg}<10'b0010011011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0010011011)) color_data = 12'b101110110011;
		if(({row_reg, col_reg}==10'b0010011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0010011101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0010100000)) color_data = 12'b111011100110;
		if(({row_reg, col_reg}==10'b0010100001)) color_data = 12'b111111110111;
		if(({row_reg, col_reg}==10'b0010100010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0010100011)) color_data = 12'b110111000110;
		if(({row_reg, col_reg}==10'b0010100100)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}>=10'b0010100101) && ({row_reg, col_reg}<10'b0010100111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0010100111) && ({row_reg, col_reg}<10'b0010101001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0010101001) && ({row_reg, col_reg}<10'b0010101011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0010101011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0010101100) && ({row_reg, col_reg}<10'b0010101111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0010101111)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0010110000)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}>=10'b0010110001) && ({row_reg, col_reg}<10'b0010111001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0010111001) && ({row_reg, col_reg}<10'b0010111011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0010111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0010111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0010111101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0011000000)) color_data = 12'b111011110110;
		if(({row_reg, col_reg}==10'b0011000001)) color_data = 12'b111111110111;
		if(({row_reg, col_reg}==10'b0011000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0011000011)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}>=10'b0011000100) && ({row_reg, col_reg}<10'b0011000110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0011000110) && ({row_reg, col_reg}<10'b0011001000)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}>=10'b0011001000) && ({row_reg, col_reg}<10'b0011001100)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0011001100)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}>=10'b0011001101) && ({row_reg, col_reg}<10'b0011001111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0011001111)) color_data = 12'b110011100101;
		if(({row_reg, col_reg}==10'b0011010000)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0011010001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0011010010) && ({row_reg, col_reg}<10'b0011011001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0011011001) && ({row_reg, col_reg}<10'b0011011011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0011011011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0011011100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b0011011101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0011100000)) color_data = 12'b111011110110;
		if(({row_reg, col_reg}==10'b0011100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0011100010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0011100011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0011100100)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0011100101)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}>=10'b0011100110) && ({row_reg, col_reg}<10'b0011101000)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}>=10'b0011101000) && ({row_reg, col_reg}<10'b0011101100)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0011101100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0011101101)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}==10'b0011101110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0011101111)) color_data = 12'b110011100101;
		if(({row_reg, col_reg}==10'b0011110000)) color_data = 12'b111110110110;
		if(({row_reg, col_reg}==10'b0011110001)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b0011110010)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0011110011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0011110100)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}>=10'b0011110101) && ({row_reg, col_reg}<10'b0011111000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0011111000) && ({row_reg, col_reg}<10'b0011111010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0011111010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0011111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0011111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0011111101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b0100000000)) color_data = 12'b111011110111;
		if(({row_reg, col_reg}==10'b0100000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0100000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0100000011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0100000100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0100000101) && ({row_reg, col_reg}<10'b0100001000)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0100001000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0100001001) && ({row_reg, col_reg}<10'b0100001110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0100001110)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0100001111)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b0100010000)) color_data = 12'b111110000101;
		if(({row_reg, col_reg}==10'b0100010001)) color_data = 12'b110001110011;
		if(({row_reg, col_reg}==10'b0100010010)) color_data = 12'b111010110101;
		if(({row_reg, col_reg}==10'b0100010011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0100010100)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0100010101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0100010110) && ({row_reg, col_reg}<10'b0100011000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0100011000) && ({row_reg, col_reg}<10'b0100011011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0100011011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0100011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0100011101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0100100000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0100100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0100100010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0100100011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0100100100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0100100101) && ({row_reg, col_reg}<10'b0100100111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0100100111)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==10'b0100101000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0100101001) && ({row_reg, col_reg}<10'b0100101011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0100101011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0100101100)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==10'b0100101101)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b0100101110)) color_data = 12'b111110110110;
		if(({row_reg, col_reg}==10'b0100101111)) color_data = 12'b111110000100;
		if(({row_reg, col_reg}==10'b0100110000)) color_data = 12'b111101000011;
		if(({row_reg, col_reg}==10'b0100110001)) color_data = 12'b110101010010;
		if(({row_reg, col_reg}==10'b0100110010)) color_data = 12'b111010100101;
		if(({row_reg, col_reg}>=10'b0100110011) && ({row_reg, col_reg}<10'b0100110101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0100110101)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0100110110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0100110111) && ({row_reg, col_reg}<10'b0100111011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0100111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0100111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0100111101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0101000000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0101000001)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==10'b0101000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b0101000011) && ({row_reg, col_reg}<10'b0101000101)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}>=10'b0101000101) && ({row_reg, col_reg}<10'b0101000111)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0101000111)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==10'b0101001000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0101001001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0101001010)) color_data = 12'b111111000101;
		if(({row_reg, col_reg}==10'b0101001011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0101001100)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b0101001101)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b0101001110)) color_data = 12'b111010000100;
		if(({row_reg, col_reg}==10'b0101001111)) color_data = 12'b111001000010;
		if(({row_reg, col_reg}==10'b0101010000)) color_data = 12'b111100100100;
		if(({row_reg, col_reg}==10'b0101010001)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b0101010010)) color_data = 12'b110110100100;
		if(({row_reg, col_reg}>=10'b0101010011) && ({row_reg, col_reg}<10'b0101010110)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}>=10'b0101010110) && ({row_reg, col_reg}<10'b0101011000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0101011000) && ({row_reg, col_reg}<10'b0101011011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0101011011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0101011100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b0101011101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0101100000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0101100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0101100010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0101100011)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}==10'b0101100100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0101100101) && ({row_reg, col_reg}<10'b0101101010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0101101010)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0101101011)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b0101101100)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b0101101101)) color_data = 12'b111010000100;
		if(({row_reg, col_reg}==10'b0101101110)) color_data = 12'b110101010010;
		if(({row_reg, col_reg}==10'b0101101111)) color_data = 12'b111001000011;
		if(({row_reg, col_reg}==10'b0101110000)) color_data = 12'b111100110101;
		if(({row_reg, col_reg}==10'b0101110001)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b0101110010)) color_data = 12'b111010100101;
		if(({row_reg, col_reg}>=10'b0101110011) && ({row_reg, col_reg}<10'b0101110110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0101110110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0101110111)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}>=10'b0101111000) && ({row_reg, col_reg}<10'b0101111010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0101111010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0101111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0101111100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b0101111101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b0110000000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0110000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0110000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b0110000011) && ({row_reg, col_reg}<10'b0110000110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0110000110) && ({row_reg, col_reg}<10'b0110001000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0110001000) && ({row_reg, col_reg}<10'b0110001010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0110001010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0110001011)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b0110001100)) color_data = 12'b111110000100;
		if(({row_reg, col_reg}==10'b0110001101)) color_data = 12'b110101000010;
		if(({row_reg, col_reg}==10'b0110001110)) color_data = 12'b110101010010;
		if(({row_reg, col_reg}==10'b0110001111)) color_data = 12'b111110010110;
		if(({row_reg, col_reg}==10'b0110010000)) color_data = 12'b111101000110;
		if(({row_reg, col_reg}==10'b0110010001)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b0110010010)) color_data = 12'b111010100101;
		if(({row_reg, col_reg}==10'b0110010011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0110010100)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0110010101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0110010110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b0110010111) && ({row_reg, col_reg}<10'b0110011010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0110011010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0110011011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0110011100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b0110011101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b0110100000)) color_data = 12'b111111100111;
		if(({row_reg, col_reg}==10'b0110100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0110100010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b0110100011) && ({row_reg, col_reg}<10'b0110100101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0110100101) && ({row_reg, col_reg}<10'b0110100111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0110100111)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}==10'b0110101000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0110101001)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==10'b0110101010)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b0110101011)) color_data = 12'b111010000100;
		if(({row_reg, col_reg}==10'b0110101100)) color_data = 12'b110101000010;
		if(({row_reg, col_reg}==10'b0110101101)) color_data = 12'b111001010011;
		if(({row_reg, col_reg}==10'b0110101110)) color_data = 12'b111110010101;
		if(({row_reg, col_reg}==10'b0110101111)) color_data = 12'b111110110110;
		if(({row_reg, col_reg}==10'b0110110000)) color_data = 12'b111101010110;
		if(({row_reg, col_reg}==10'b0110110001)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b0110110010)) color_data = 12'b111010100101;
		if(({row_reg, col_reg}==10'b0110110011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0110110100)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0110110101)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0110110110)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0110110111)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b0110111000) && ({row_reg, col_reg}<10'b0110111010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0110111010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0110111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b0110111100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b0110111101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b0111000000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0111000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0111000010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b0111000011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b0111000100) && ({row_reg, col_reg}<10'b0111000110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0111000110)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}==10'b0111000111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0111001000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0111001001)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b0111001010)) color_data = 12'b111010100110;
		if(({row_reg, col_reg}>=10'b0111001011) && ({row_reg, col_reg}<10'b0111001101)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b0111001101)) color_data = 12'b111110010110;
		if(({row_reg, col_reg}==10'b0111001110)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b0111001111)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}==10'b0111010000)) color_data = 12'b111101000101;
		if(({row_reg, col_reg}==10'b0111010001)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b0111010010)) color_data = 12'b111010100100;
		if(({row_reg, col_reg}==10'b0111010011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}>=10'b0111010100) && ({row_reg, col_reg}<10'b0111010110)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b0111010110)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}>=10'b0111010111) && ({row_reg, col_reg}<10'b0111011001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0111011001)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0111011010)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}==10'b0111011011)) color_data = 12'b110010110011;
		if(({row_reg, col_reg}==10'b0111011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0111011101)) color_data = 12'b100110100011;
		if(({row_reg, col_reg}==10'b0111100000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b0111100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b0111100010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b0111100011)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}==10'b0111100100)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0111100101)) color_data = 12'b111011000100;
		if(({row_reg, col_reg}==10'b0111100110)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0111100111)) color_data = 12'b110011100100;
		if(({row_reg, col_reg}==10'b0111101000)) color_data = 12'b110011010100;
		if(({row_reg, col_reg}==10'b0111101001)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b0111101010)) color_data = 12'b111110000101;
		if(({row_reg, col_reg}==10'b0111101011)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b0111101100)) color_data = 12'b110101010100;
		if(({row_reg, col_reg}==10'b0111101101)) color_data = 12'b111010010101;
		if(({row_reg, col_reg}==10'b0111101110)) color_data = 12'b110010010011;
		if(({row_reg, col_reg}==10'b0111101111)) color_data = 12'b101110100010;
		if(({row_reg, col_reg}==10'b0111110000)) color_data = 12'b111101000101;
		if(({row_reg, col_reg}==10'b0111110001)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b0111110010)) color_data = 12'b110110000011;
		if(({row_reg, col_reg}==10'b0111110011)) color_data = 12'b110110110011;
		if(({row_reg, col_reg}>=10'b0111110100) && ({row_reg, col_reg}<10'b0111110110)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b0111110110)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b0111110111)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b0111111000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b0111111001)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b0111111010)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}==10'b0111111011)) color_data = 12'b110010110011;
		if(({row_reg, col_reg}==10'b0111111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b0111111101)) color_data = 12'b100110100011;
		if(({row_reg, col_reg}==10'b1000000000)) color_data = 12'b111111100111;
		if(({row_reg, col_reg}==10'b1000000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1000000010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1000000011) && ({row_reg, col_reg}<10'b1000000111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b1000000111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1000001000)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1000001001)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b1000001010)) color_data = 12'b111010010101;
		if(({row_reg, col_reg}==10'b1000001011)) color_data = 12'b110001010010;
		if(({row_reg, col_reg}==10'b1000001100)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b1000001101)) color_data = 12'b111000110011;
		if(({row_reg, col_reg}>=10'b1000001110) && ({row_reg, col_reg}<10'b1000010000)) color_data = 12'b111100110011;
		if(({row_reg, col_reg}>=10'b1000010000) && ({row_reg, col_reg}<10'b1000010010)) color_data = 12'b111100110100;
		if(({row_reg, col_reg}==10'b1000010010)) color_data = 12'b111000110010;
		if(({row_reg, col_reg}==10'b1000010011)) color_data = 12'b110101010010;
		if(({row_reg, col_reg}==10'b1000010100)) color_data = 12'b111110110110;
		if(({row_reg, col_reg}>=10'b1000010101) && ({row_reg, col_reg}<10'b1000011000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1000011000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1000011001)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1000011010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1000011011)) color_data = 12'b101110110100;
		if(({row_reg, col_reg}==10'b1000011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1000011101)) color_data = 12'b100110100011;
		if(({row_reg, col_reg}==10'b1000100000)) color_data = 12'b111111100111;
		if(({row_reg, col_reg}==10'b1000100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1000100010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b1000100011) && ({row_reg, col_reg}<10'b1000100101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1000100101) && ({row_reg, col_reg}<10'b1000100111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b1000100111)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1000101000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1000101001)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b1000101010)) color_data = 12'b111010110101;
		if(({row_reg, col_reg}==10'b1000101011)) color_data = 12'b110110000100;
		if(({row_reg, col_reg}==10'b1000101100)) color_data = 12'b110101110100;
		if(({row_reg, col_reg}==10'b1000101101)) color_data = 12'b111001110100;
		if(({row_reg, col_reg}>=10'b1000101110) && ({row_reg, col_reg}<10'b1000110000)) color_data = 12'b111001100100;
		if(({row_reg, col_reg}==10'b1000110000)) color_data = 12'b111001000100;
		if(({row_reg, col_reg}==10'b1000110001)) color_data = 12'b111001000011;
		if(({row_reg, col_reg}==10'b1000110010)) color_data = 12'b111001100100;
		if(({row_reg, col_reg}==10'b1000110011)) color_data = 12'b110110000100;
		if(({row_reg, col_reg}==10'b1000110100)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}>=10'b1000110101) && ({row_reg, col_reg}<10'b1000110111)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==10'b1000110111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}>=10'b1000111000) && ({row_reg, col_reg}<10'b1000111011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1000111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b1000111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1000111101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b1001000000)) color_data = 12'b111111101000;
		if(({row_reg, col_reg}==10'b1001000001)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==10'b1001000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b1001000011) && ({row_reg, col_reg}<10'b1001000101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1001000101) && ({row_reg, col_reg}<10'b1001001000)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}>=10'b1001001000) && ({row_reg, col_reg}<10'b1001001010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1001001010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1001001011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1001001100)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}>=10'b1001001101) && ({row_reg, col_reg}<10'b1001010000)) color_data = 12'b111111000110;
		if(({row_reg, col_reg}==10'b1001010000)) color_data = 12'b111101010100;
		if(({row_reg, col_reg}==10'b1001010001)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b1001010010)) color_data = 12'b111010010110;
		if(({row_reg, col_reg}==10'b1001010011)) color_data = 12'b111011000111;
		if(({row_reg, col_reg}==10'b1001010100)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b1001010101) && ({row_reg, col_reg}<10'b1001011011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1001011011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b1001011100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b1001011101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b1001100000)) color_data = 12'b111011101000;
		if(({row_reg, col_reg}==10'b1001100001)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==10'b1001100010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b1001100011) && ({row_reg, col_reg}<10'b1001101101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1001101101) && ({row_reg, col_reg}<10'b1001110000)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b1001110000)) color_data = 12'b111101010100;
		if(({row_reg, col_reg}==10'b1001110001)) color_data = 12'b110001000010;
		if(({row_reg, col_reg}==10'b1001110010)) color_data = 12'b111010100110;
		if(({row_reg, col_reg}==10'b1001110011)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b1001110100)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}==10'b1001110101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1001110110) && ({row_reg, col_reg}<10'b1001111000)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}>=10'b1001111000) && ({row_reg, col_reg}<10'b1001111011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1001111011)) color_data = 12'b101110110100;
		if(({row_reg, col_reg}==10'b1001111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1001111101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1010000000)) color_data = 12'b111011101000;
		if(({row_reg, col_reg}==10'b1010000001)) color_data = 12'b111111111001;
		if(({row_reg, col_reg}==10'b1010000010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b1010000011) && ({row_reg, col_reg}<10'b1010000110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1010000110) && ({row_reg, col_reg}<10'b1010001001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010001001)) color_data = 12'b110111000101;
		if(({row_reg, col_reg}>=10'b1010001010) && ({row_reg, col_reg}<10'b1010001100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010001100)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1010001101) && ({row_reg, col_reg}<10'b1010010000)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b1010010000)) color_data = 12'b111101010011;
		if(({row_reg, col_reg}==10'b1010010001)) color_data = 12'b110001000001;
		if(({row_reg, col_reg}==10'b1010010010)) color_data = 12'b111010100101;
		if(({row_reg, col_reg}==10'b1010010011)) color_data = 12'b111011000110;
		if(({row_reg, col_reg}==10'b1010010100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010010101)) color_data = 12'b111111010101;
		if(({row_reg, col_reg}==10'b1010010110)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1010010111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1010011000) && ({row_reg, col_reg}<10'b1010011011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1010011011)) color_data = 12'b101110110100;
		if(({row_reg, col_reg}==10'b1010011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1010011101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1010100000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b1010100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1010100010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b1010100011) && ({row_reg, col_reg}<10'b1010100101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1010100101) && ({row_reg, col_reg}<10'b1010100111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1010100111) && ({row_reg, col_reg}<10'b1010101001)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1010101001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010101010)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1010101011)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010101100)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}>=10'b1010101101) && ({row_reg, col_reg}<10'b1010101111)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010101111)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}==10'b1010110000)) color_data = 12'b111101110011;
		if(({row_reg, col_reg}==10'b1010110001)) color_data = 12'b110001110010;
		if(({row_reg, col_reg}==10'b1010110010)) color_data = 12'b111010110101;
		if(({row_reg, col_reg}==10'b1010110011)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1010110100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1010110101)) color_data = 12'b111111000101;
		if(({row_reg, col_reg}==10'b1010110110)) color_data = 12'b111011000100;
		if(({row_reg, col_reg}==10'b1010110111)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}>=10'b1010111000) && ({row_reg, col_reg}<10'b1010111011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1010111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b1010111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1010111101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1011000000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b1011000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}>=10'b1011000010) && ({row_reg, col_reg}<10'b1011000110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1011000110) && ({row_reg, col_reg}<10'b1011001000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1011001000) && ({row_reg, col_reg}<10'b1011001101)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}>=10'b1011001101) && ({row_reg, col_reg}<10'b1011010000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1011010000)) color_data = 12'b111110110110;
		if(({row_reg, col_reg}==10'b1011010001)) color_data = 12'b111010110101;
		if(({row_reg, col_reg}==10'b1011010010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b1011010011)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1011010100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1011010101) && ({row_reg, col_reg}<10'b1011010111)) color_data = 12'b111011010100;
		if(({row_reg, col_reg}>=10'b1011010111) && ({row_reg, col_reg}<10'b1011011010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1011011010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1011011011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b1011011100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b1011011101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b1011100000)) color_data = 12'b111111100111;
		if(({row_reg, col_reg}==10'b1011100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1011100010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1011100011) && ({row_reg, col_reg}<10'b1011101001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1011101001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1011101010) && ({row_reg, col_reg}<10'b1011110000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1011110000)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}>=10'b1011110001) && ({row_reg, col_reg}<10'b1011111010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1011111010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1011111011)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b1011111100)) color_data = 12'b101010010010;

		if(({row_reg, col_reg}==10'b1011111101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b1100000000)) color_data = 12'b111111100111;
		if(({row_reg, col_reg}==10'b1100000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1100000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b1100000011) && ({row_reg, col_reg}<10'b1100010000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1100010000)) color_data = 12'b110011010101;
		if(({row_reg, col_reg}==10'b1100010001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1100010010) && ({row_reg, col_reg}<10'b1100010100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1100010100) && ({row_reg, col_reg}<10'b1100011010)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1100011010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b1100011011)) color_data = 12'b101111000100;
		if(({row_reg, col_reg}==10'b1100011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1100011101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1100100000)) color_data = 12'b111111100111;
		if(({row_reg, col_reg}==10'b1100100001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1100100010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}>=10'b1100100011) && ({row_reg, col_reg}<10'b1100101000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1100101000) && ({row_reg, col_reg}<10'b1100101100)) color_data = 12'b110111010100;
		if(({row_reg, col_reg}>=10'b1100101100) && ({row_reg, col_reg}<10'b1100110001)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}==10'b1100110001)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1100110010) && ({row_reg, col_reg}<10'b1100110100)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1100110100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1100110101) && ({row_reg, col_reg}<10'b1100111000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1100111000) && ({row_reg, col_reg}<10'b1100111010)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1100111010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b1100111011)) color_data = 12'b101111000100;
		if(({row_reg, col_reg}==10'b1100111100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1100111101)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1101000000)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b1101000001)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1101000010)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b1101000011)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b1101000100)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b1101000101)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1101000110) && ({row_reg, col_reg}<10'b1101010000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1101010000)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1101010001) && ({row_reg, col_reg}<10'b1101010100)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}>=10'b1101010100) && ({row_reg, col_reg}<10'b1101010110)) color_data = 12'b110111010101;
		if(({row_reg, col_reg}>=10'b1101010110) && ({row_reg, col_reg}<10'b1101011000)) color_data = 12'b111011010101;
		if(({row_reg, col_reg}==10'b1101011000)) color_data = 12'b111011000101;
		if(({row_reg, col_reg}==10'b1101011001)) color_data = 12'b111011010110;
		if(({row_reg, col_reg}==10'b1101011010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b1101011011)) color_data = 12'b101110110100;
		if(({row_reg, col_reg}==10'b1101011100)) color_data = 12'b100110010010;

		if(({row_reg, col_reg}==10'b1101011101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}>=10'b1101100000) && ({row_reg, col_reg}<10'b1101100010)) color_data = 12'b111111111000;
		if(({row_reg, col_reg}==10'b1101100010)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b1101100011)) color_data = 12'b101110100100;
		if(({row_reg, col_reg}>=10'b1101100100) && ({row_reg, col_reg}<10'b1101100110)) color_data = 12'b101110100011;
		if(({row_reg, col_reg}==10'b1101100110)) color_data = 12'b101110110011;
		if(({row_reg, col_reg}>=10'b1101100111) && ({row_reg, col_reg}<10'b1101101101)) color_data = 12'b101110100011;
		if(({row_reg, col_reg}>=10'b1101101101) && ({row_reg, col_reg}<10'b1101110000)) color_data = 12'b101110100100;
		if(({row_reg, col_reg}>=10'b1101110000) && ({row_reg, col_reg}<10'b1101110100)) color_data = 12'b101110110011;
		if(({row_reg, col_reg}==10'b1101110100)) color_data = 12'b101010110011;
		if(({row_reg, col_reg}>=10'b1101110101) && ({row_reg, col_reg}<10'b1101110111)) color_data = 12'b101110110011;
		if(({row_reg, col_reg}>=10'b1101110111) && ({row_reg, col_reg}<10'b1101111001)) color_data = 12'b110010100011;
		if(({row_reg, col_reg}==10'b1101111001)) color_data = 12'b101110100011;
		if(({row_reg, col_reg}==10'b1101111010)) color_data = 12'b101110110100;
		if(({row_reg, col_reg}==10'b1101111011)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1101111100)) color_data = 12'b100110000010;

		if(({row_reg, col_reg}==10'b1101111101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}==10'b1110000000)) color_data = 12'b110111010110;
		if(({row_reg, col_reg}==10'b1110000001)) color_data = 12'b111011100111;
		if(({row_reg, col_reg}==10'b1110000010)) color_data = 12'b101110110100;
		if(({row_reg, col_reg}>=10'b1110000011) && ({row_reg, col_reg}<10'b1110000110)) color_data = 12'b100110010010;
		if(({row_reg, col_reg}>=10'b1110000110) && ({row_reg, col_reg}<10'b1110001100)) color_data = 12'b101010010010;
		if(({row_reg, col_reg}==10'b1110001100)) color_data = 12'b100110010010;
		if(({row_reg, col_reg}>=10'b1110001101) && ({row_reg, col_reg}<10'b1110010000)) color_data = 12'b100110010011;
		if(({row_reg, col_reg}>=10'b1110010000) && ({row_reg, col_reg}<10'b1110010111)) color_data = 12'b100110010010;
		if(({row_reg, col_reg}>=10'b1110010111) && ({row_reg, col_reg}<10'b1110011001)) color_data = 12'b101010010010;
		if(({row_reg, col_reg}>=10'b1110011001) && ({row_reg, col_reg}<10'b1110011100)) color_data = 12'b100110010010;
		if(({row_reg, col_reg}==10'b1110011100)) color_data = 12'b100010000010;

		if(({row_reg, col_reg}==10'b1110011101)) color_data = 12'b100110000010;
		if(({row_reg, col_reg}==10'b1110100000)) color_data = 12'b110010110100;
		if(({row_reg, col_reg}==10'b1110100001)) color_data = 12'b110011000100;
		if(({row_reg, col_reg}==10'b1110100010)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1110100011)) color_data = 12'b101010010010;
		if(({row_reg, col_reg}==10'b1110100100)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1110100101)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}>=10'b1110100110) && ({row_reg, col_reg}<10'b1110101000)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}>=10'b1110101000) && ({row_reg, col_reg}<10'b1110101010)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}>=10'b1110101010) && ({row_reg, col_reg}<10'b1110110000)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1110110000)) color_data = 12'b101010010011;
		if(({row_reg, col_reg}>=10'b1110110001) && ({row_reg, col_reg}<10'b1110110011)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1110110011)) color_data = 12'b100110100011;
		if(({row_reg, col_reg}>=10'b1110110100) && ({row_reg, col_reg}<10'b1110111011)) color_data = 12'b101010100011;
		if(({row_reg, col_reg}==10'b1110111011)) color_data = 12'b100110010011;
		if(({row_reg, col_reg}==10'b1110111100)) color_data = 12'b100010000010;

		if(({row_reg, col_reg}>=10'b1110111101) && ({row_reg, col_reg}<=10'b1110111101)) color_data = 12'b011101110001;
	end
endmodule