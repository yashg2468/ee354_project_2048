module tile_rom_1024
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==10'b0000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==10'b0000000001)) color_data = 12'b111111001101;
		if(({row_reg, col_reg}==10'b0000000010)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b0000000011)) color_data = 12'b111110001011;
		if(({row_reg, col_reg}==10'b0000000100)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b0000000101)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}>=10'b0000000110) && ({row_reg, col_reg}<10'b0000001001)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}>=10'b0000001001) && ({row_reg, col_reg}<10'b0000001011)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0000001011)) color_data = 12'b111110001011;
		if(({row_reg, col_reg}>=10'b0000001100) && ({row_reg, col_reg}<10'b0000001110)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}>=10'b0000001110) && ({row_reg, col_reg}<10'b0000010000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0000010000)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}==10'b0000010001)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}>=10'b0000010010) && ({row_reg, col_reg}<10'b0000010111)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0000010111)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b0000011000)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}==10'b0000011001)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b0000011010)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0000011011)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}==10'b0000011100)) color_data = 12'b111001000111;

		if(({row_reg, col_reg}==10'b0000011101)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}>=10'b0000100000) && ({row_reg, col_reg}<10'b0000100010)) color_data = 12'b111111001101;
		if(({row_reg, col_reg}==10'b0000100010)) color_data = 12'b111110101100;
		if(({row_reg, col_reg}>=10'b0000100011) && ({row_reg, col_reg}<10'b0000111011)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0000111011)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b0000111100)) color_data = 12'b110000110110;

		if(({row_reg, col_reg}==10'b0000111101)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b0001000000)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}>=10'b0001000001) && ({row_reg, col_reg}<10'b0001000011)) color_data = 12'b111110101100;
		if(({row_reg, col_reg}>=10'b0001000011) && ({row_reg, col_reg}<10'b0001000101)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}==10'b0001000101)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}>=10'b0001000110) && ({row_reg, col_reg}<10'b0001001000)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}==10'b0001001000)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}>=10'b0001001001) && ({row_reg, col_reg}<10'b0001001110)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}>=10'b0001001110) && ({row_reg, col_reg}<10'b0001010000)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0001010000)) color_data = 12'b111101101010;
		if(({row_reg, col_reg}>=10'b0001010001) && ({row_reg, col_reg}<10'b0001010101)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}>=10'b0001010101) && ({row_reg, col_reg}<10'b0001011010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0001011010)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}==10'b0001011011)) color_data = 12'b110000110110;

		if(({row_reg, col_reg}>=10'b0001011100) && ({row_reg, col_reg}<10'b0001100000)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}>=10'b0001100000) && ({row_reg, col_reg}<10'b0001100010)) color_data = 12'b111110001011;
		if(({row_reg, col_reg}==10'b0001100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0001100011)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}>=10'b0001100100) && ({row_reg, col_reg}<10'b0001100110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0001100110)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b0001100111) && ({row_reg, col_reg}<10'b0001101010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b0001101010) && ({row_reg, col_reg}<10'b0001101100)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b0001101100) && ({row_reg, col_reg}<10'b0001101111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0001101111)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0001110000)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0001110001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0001110010)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b0001110011) && ({row_reg, col_reg}<10'b0001110111)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}>=10'b0001110111) && ({row_reg, col_reg}<10'b0001111010)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0001111010)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b0001111011)) color_data = 12'b101000010100;

		if(({row_reg, col_reg}>=10'b0001111100) && ({row_reg, col_reg}<10'b0010000000)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}>=10'b0010000000) && ({row_reg, col_reg}<10'b0010000010)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0010000010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b0010000011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b0010000100) && ({row_reg, col_reg}<10'b0010000110)) color_data = 12'b111101000111;
		if(({row_reg, col_reg}>=10'b0010000110) && ({row_reg, col_reg}<10'b0010001001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010001001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b0010001010) && ({row_reg, col_reg}<10'b0010011000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010011000)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0010011001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010011010)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0010011011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b0010011100)) color_data = 12'b101000100101;

		if(({row_reg, col_reg}==10'b0010011101)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==10'b0010100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0010100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0010100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}>=10'b0010100011) && ({row_reg, col_reg}<10'b0010100110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010100110)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b0010100111) && ({row_reg, col_reg}<10'b0010101001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010101001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b0010101010) && ({row_reg, col_reg}<10'b0010101100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010101100)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}>=10'b0010101101) && ({row_reg, col_reg}<10'b0010101111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0010101111)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}==10'b0010110000)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}>=10'b0010110001) && ({row_reg, col_reg}<10'b0010111001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b0010111001) && ({row_reg, col_reg}<10'b0010111011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0010111011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b0010111100)) color_data = 12'b101000100101;

		if(({row_reg, col_reg}==10'b0010111101)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b0011000000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0011000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0011000010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0011000011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b0011000100) && ({row_reg, col_reg}<10'b0011001100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b0011001100) && ({row_reg, col_reg}<10'b0011001110)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0011001110)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0011001111)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0011010000)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}>=10'b0011010001) && ({row_reg, col_reg}<10'b0011010100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0011010100)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0011010101)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0011010110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0011010111)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0011011000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0011011001)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b0011011010)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0011011011)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0011011100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b0011011101)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}>=10'b0011100000) && ({row_reg, col_reg}<10'b0011100010)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0011100010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b0011100011)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0011100100)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}>=10'b0011100101) && ({row_reg, col_reg}<10'b0011110010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0011110010)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0011110011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0011110100)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0011110101)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}>=10'b0011110110) && ({row_reg, col_reg}<10'b0011111001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b0011111001) && ({row_reg, col_reg}<10'b0011111011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0011111011)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0011111100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b0011111101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b0100000000)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}==10'b0100000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0100000010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0100000011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0100000100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100000101)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0100000110)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b0100000111) && ({row_reg, col_reg}<10'b0100001001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100001001)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b0100001010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}==10'b0100001011)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}>=10'b0100001100) && ({row_reg, col_reg}<10'b0100001110)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b0100001110)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0100001111)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}>=10'b0100010000) && ({row_reg, col_reg}<10'b0100010100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100010100)) color_data = 12'b111101000111;
		if(({row_reg, col_reg}>=10'b0100010101) && ({row_reg, col_reg}<10'b0100010111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b0100010111) && ({row_reg, col_reg}<10'b0100011010)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0100011010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100011011)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==10'b0100011100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b0100011101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b0100100000)) color_data = 12'b111010011011;
		if(({row_reg, col_reg}==10'b0100100001)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0100100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0100100011)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b0100100100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100100101)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0100100110)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b0100100111)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}>=10'b0100101000) && ({row_reg, col_reg}<10'b0100101011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100101011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b0100101100)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==10'b0100101101)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0100101110)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0100101111)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0100110000)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0100110001)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b0100110010)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==10'b0100110011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100110100)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b0100110101)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0100110110)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0100110111)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0100111000)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0100111001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0100111010)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b0100111011)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0100111100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b0100111101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b0101000000)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b0101000001)) color_data = 12'b111110011100;
		if(({row_reg, col_reg}==10'b0101000010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}>=10'b0101000011) && ({row_reg, col_reg}<10'b0101000101)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b0101000101)) color_data = 12'b110001000111;
		if(({row_reg, col_reg}==10'b0101000110)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==10'b0101000111)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0101001000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0101001001)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0101001010)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}>=10'b0101001011) && ({row_reg, col_reg}<10'b0101001101)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==10'b0101001101)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0101001110)) color_data = 12'b101001000110;
		if(({row_reg, col_reg}==10'b0101001111)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b0101010000)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==10'b0101010001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==10'b0101010010)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==10'b0101010011)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==10'b0101010100)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b0101010101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0101010110)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==10'b0101010111)) color_data = 12'b010000000001;
		if(({row_reg, col_reg}==10'b0101011000)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}>=10'b0101011001) && ({row_reg, col_reg}<10'b0101011011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0101011011)) color_data = 12'b101100100101;

		if(({row_reg, col_reg}>=10'b0101011100) && ({row_reg, col_reg}<10'b0101100000)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b0101100000)) color_data = 12'b111110001011;
		if(({row_reg, col_reg}==10'b0101100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0101100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b0101100011)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==10'b0101100100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0101100101)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b0101100110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==10'b0101100111)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0101101000)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b0101101001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0101101010)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b0101101011)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==10'b0101101100)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==10'b0101101101)) color_data = 12'b010000000001;
		if(({row_reg, col_reg}==10'b0101101110)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==10'b0101101111)) color_data = 12'b011000010010;
		if(({row_reg, col_reg}==10'b0101110000)) color_data = 12'b100000100011;
		if(({row_reg, col_reg}==10'b0101110001)) color_data = 12'b100001010101;
		if(({row_reg, col_reg}==10'b0101110010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==10'b0101110011)) color_data = 12'b011100010010;
		if(({row_reg, col_reg}==10'b0101110100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0101110101)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b0101110110)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==10'b0101110111)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==10'b0101111000)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==10'b0101111001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0101111010)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b0101111011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b0101111100)) color_data = 12'b100100100100;

		if(({row_reg, col_reg}==10'b0101111101)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b0110000000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0110000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0110000010)) color_data = 12'b111001111001;
		if(({row_reg, col_reg}==10'b0110000011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0110000100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0110000101)) color_data = 12'b011100000001;
		if(({row_reg, col_reg}==10'b0110000110)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==10'b0110000111)) color_data = 12'b011000000010;
		if(({row_reg, col_reg}>=10'b0110001000) && ({row_reg, col_reg}<10'b0110001010)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0110001010)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==10'b0110001011)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==10'b0110001100)) color_data = 12'b101101010111;
		if(({row_reg, col_reg}==10'b0110001101)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b0110001110)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b0110001111)) color_data = 12'b100100110101;
		if(({row_reg, col_reg}==10'b0110010000)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0110010001)) color_data = 12'b101101010111;
		if(({row_reg, col_reg}==10'b0110010010)) color_data = 12'b011100110100;
		if(({row_reg, col_reg}==10'b0110010011)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==10'b0110010100)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b0110010101)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b0110010110)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==10'b0110010111)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0110011000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0110011001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b0110011010)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b0110011011)) color_data = 12'b101000100101;

		if(({row_reg, col_reg}>=10'b0110011100) && ({row_reg, col_reg}<10'b0110100000)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b0110100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0110100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0110100010)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0110100011)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0110100100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0110100101)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0110100110)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==10'b0110100111)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b0110101000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0110101001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0110101010)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==10'b0110101011)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==10'b0110101100)) color_data = 12'b110001000111;
		if(({row_reg, col_reg}==10'b0110101101)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==10'b0110101110)) color_data = 12'b101000000011;
		if(({row_reg, col_reg}==10'b0110101111)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b0110110000)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b0110110001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0110110010)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==10'b0110110011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b0110110100)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b0110110101)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0110110110)) color_data = 12'b011100110100;
		if(({row_reg, col_reg}==10'b0110110111)) color_data = 12'b011000000010;
		if(({row_reg, col_reg}==10'b0110111000)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b0110111001)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b0110111010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0110111011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b0110111100)) color_data = 12'b100100110101;

		if(({row_reg, col_reg}==10'b0110111101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b0111000000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0111000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b0111000010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b0111000011)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0111000100)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0111000101)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0111000110)) color_data = 12'b101101000101;
		if(({row_reg, col_reg}==10'b0111000111)) color_data = 12'b011100000001;
		if(({row_reg, col_reg}==10'b0111001000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0111001001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0111001010)) color_data = 12'b100000000001;
		if(({row_reg, col_reg}==10'b0111001011)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==10'b0111001100)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}>=10'b0111001101) && ({row_reg, col_reg}<10'b0111001111)) color_data = 12'b101000000011;
		if(({row_reg, col_reg}==10'b0111001111)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0111010000)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0111010001)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b0111010010)) color_data = 12'b010100000000;
		if(({row_reg, col_reg}==10'b0111010011)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==10'b0111010100)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==10'b0111010101)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==10'b0111010110)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}==10'b0111010111)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0111011000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0111011001)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b0111011010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0111011011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b0111011100)) color_data = 12'b101000110101;

		if(({row_reg, col_reg}==10'b0111011101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b0111100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b0111100001)) color_data = 12'b111110001011;
		if(({row_reg, col_reg}==10'b0111100010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}>=10'b0111100011) && ({row_reg, col_reg}<10'b0111100101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b0111100101)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b0111100110)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==10'b0111100111)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b0111101000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b0111101001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b0111101010)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==10'b0111101011)) color_data = 12'b101001000101;
		if(({row_reg, col_reg}==10'b0111101100)) color_data = 12'b110001010111;
		if(({row_reg, col_reg}==10'b0111101101)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b0111101110)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b0111101111)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0111110000)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==10'b0111110001)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b0111110010)) color_data = 12'b011100000011;
		if(({row_reg, col_reg}==10'b0111110011)) color_data = 12'b101001010110;
		if(({row_reg, col_reg}==10'b0111110100)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==10'b0111110101)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==10'b0111110110)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==10'b0111110111)) color_data = 12'b010000000000;
		if(({row_reg, col_reg}==10'b0111111000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b0111111001)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b0111111010)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b0111111011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b0111111100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b0111111101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1000000000)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}==10'b1000000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1000000010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b1000000011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1000000100)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1000000101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1000000110)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b1000000111)) color_data = 12'b011100000001;
		if(({row_reg, col_reg}>=10'b1000001000) && ({row_reg, col_reg}<10'b1000001010)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1000001010)) color_data = 12'b011100000001;
		if(({row_reg, col_reg}==10'b1000001011)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b1000001100)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1000001101)) color_data = 12'b101100000100;
		if(({row_reg, col_reg}==10'b1000001110)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b1000001111)) color_data = 12'b101001010111;
		if(({row_reg, col_reg}==10'b1000010000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==10'b1000010001)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b1000010010)) color_data = 12'b110100100110;
		if(({row_reg, col_reg}==10'b1000010011)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1000010100)) color_data = 12'b101100000011;
		if(({row_reg, col_reg}==10'b1000010101)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==10'b1000010110)) color_data = 12'b010000010001;
		if(({row_reg, col_reg}==10'b1000010111)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==10'b1000011000)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b1000011001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1000011010)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}>=10'b1000011011) && ({row_reg, col_reg}<10'b1000011101)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b1000011101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1000100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b1000100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1000100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}>=10'b1000100011) && ({row_reg, col_reg}<10'b1000100101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1000100101)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b1000100110)) color_data = 12'b100101010110;
		if(({row_reg, col_reg}==10'b1000100111)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==10'b1000101000)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==10'b1000101001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b1000101010)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b1000101011)) color_data = 12'b100100110101;
		if(({row_reg, col_reg}==10'b1000101100)) color_data = 12'b101101010111;
		if(({row_reg, col_reg}==10'b1000101101)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==10'b1000101110)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b1000101111)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==10'b1000110000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==10'b1000110001)) color_data = 12'b100001010101;
		if(({row_reg, col_reg}==10'b1000110010)) color_data = 12'b110001010111;
		if(({row_reg, col_reg}==10'b1000110011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1000110100)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b1000110101)) color_data = 12'b101101000110;
		if(({row_reg, col_reg}==10'b1000110110)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==10'b1000110111)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b1000111000)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b1000111001)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b1000111010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1000111011)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==10'b1000111100)) color_data = 12'b101100100101;

		if(({row_reg, col_reg}==10'b1000111101)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1001000000)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}==10'b1001000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1001000010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b1001000011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1001000100)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b1001000101)) color_data = 12'b100000110100;
		if(({row_reg, col_reg}==10'b1001000110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==10'b1001000111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==10'b1001001000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b1001001001)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b1001001010)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==10'b1001001011)) color_data = 12'b010000000001;
		if(({row_reg, col_reg}==10'b1001001100)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==10'b1001001101)) color_data = 12'b001100000000;
		if(({row_reg, col_reg}==10'b1001001110)) color_data = 12'b100100110101;
		if(({row_reg, col_reg}==10'b1001001111)) color_data = 12'b011000000010;
		if(({row_reg, col_reg}==10'b1001010000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==10'b1001010001)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==10'b1001010010)) color_data = 12'b011000010010;
		if(({row_reg, col_reg}==10'b1001010011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1001010100)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b1001010101)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b1001010110)) color_data = 12'b101001000101;
		if(({row_reg, col_reg}==10'b1001010111)) color_data = 12'b011000000010;
		if(({row_reg, col_reg}==10'b1001011000)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b1001011001)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1001011010)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b1001011011)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==10'b1001011100)) color_data = 12'b101100100101;

		if(({row_reg, col_reg}==10'b1001011101)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==10'b1001100000)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}==10'b1001100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1001100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b1001100011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1001100100)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b1001100101)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==10'b1001100110)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b1001100111)) color_data = 12'b010100000010;
		if(({row_reg, col_reg}==10'b1001101000)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==10'b1001101001)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b1001101010)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==10'b1001101011)) color_data = 12'b011000000010;
		if(({row_reg, col_reg}==10'b1001101100)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b1001101101)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b1001101110)) color_data = 12'b110001000110;
		if(({row_reg, col_reg}==10'b1001101111)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b1001110000)) color_data = 12'b010100000010;
		if(({row_reg, col_reg}==10'b1001110001)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==10'b1001110010)) color_data = 12'b011000000001;
		if(({row_reg, col_reg}==10'b1001110011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1001110100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1001110101)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b1001110110)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==10'b1001110111)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==10'b1001111000)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1001111001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1001111010)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1001111011)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==10'b1001111100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b1001111101)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==10'b1010000000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b1010000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1010000010)) color_data = 12'b111101111010;
		if(({row_reg, col_reg}==10'b1010000011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010000100)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1010000101)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}>=10'b1010000110) && ({row_reg, col_reg}<10'b1010001000)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b1010001000)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}==10'b1010001001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010001010)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1010001011)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}>=10'b1010001100) && ({row_reg, col_reg}<10'b1010001111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010001111)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b1010010000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010010001)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b1010010010)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}>=10'b1010010011) && ({row_reg, col_reg}<10'b1010010101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010010101)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}==10'b1010010110)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}>=10'b1010010111) && ({row_reg, col_reg}<10'b1010011010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010011010)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1010011011)) color_data = 12'b101100100100;

		if(({row_reg, col_reg}>=10'b1010011100) && ({row_reg, col_reg}<10'b1010100000)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1010100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b1010100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1010100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b1010100011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1010100100)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b1010100101)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1010100110)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b1010100111)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=10'b1010101000) && ({row_reg, col_reg}<10'b1010101010)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1010101010) && ({row_reg, col_reg}<10'b1010101100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010101100)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b1010101101)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1010101110)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1010101111)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1010110000)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b1010110001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1010110010)) color_data = 12'b111100100110;
		if(({row_reg, col_reg}==10'b1010110011)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1010110100)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}>=10'b1010110101) && ({row_reg, col_reg}<10'b1010111000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1010111000)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b1010111001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1010111010)) color_data = 12'b110001000110;

		if(({row_reg, col_reg}>=10'b1010111011) && ({row_reg, col_reg}<10'b1011000000)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1011000000)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b1011000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1011000010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b1011000011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b1011000100) && ({row_reg, col_reg}<10'b1011000110)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1011000110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011000111)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}>=10'b1011001000) && ({row_reg, col_reg}<10'b1011001011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011001011)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1011001100) && ({row_reg, col_reg}<10'b1011001111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b1011001111) && ({row_reg, col_reg}<10'b1011010001)) color_data = 12'b111100110111;
		if(({row_reg, col_reg}==10'b1011010001)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1011010010)) color_data = 12'b111000100110;
		if(({row_reg, col_reg}>=10'b1011010011) && ({row_reg, col_reg}<10'b1011010110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011010110)) color_data = 12'b111101000111;
		if(({row_reg, col_reg}>=10'b1011010111) && ({row_reg, col_reg}<10'b1011011001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011011001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1011011010)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b1011011011)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b1011011100)) color_data = 12'b101100100100;

		if(({row_reg, col_reg}==10'b1011011101)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==10'b1011100000)) color_data = 12'b111010011010;
		if(({row_reg, col_reg}==10'b1011100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1011100010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b1011100011)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}>=10'b1011100100) && ({row_reg, col_reg}<10'b1011100110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011100110)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}==10'b1011100111)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b1011101000) && ({row_reg, col_reg}<10'b1011101011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011101011)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1011101100)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b1011101101)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b1011101110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011101111)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1011110000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011110001)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1011110010)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}==10'b1011110011)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}==10'b1011110100)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b1011110101) && ({row_reg, col_reg}<10'b1011110111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011110111)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1011111000) && ({row_reg, col_reg}<10'b1011111010)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1011111010)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}>=10'b1011111011) && ({row_reg, col_reg}<10'b1011111101)) color_data = 12'b101100100100;

		if(({row_reg, col_reg}==10'b1011111101)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1100000000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b1100000001)) color_data = 12'b111110001011;
		if(({row_reg, col_reg}==10'b1100000010)) color_data = 12'b111101101001;
		if(({row_reg, col_reg}==10'b1100000011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100000100)) color_data = 12'b111000110111;
		if(({row_reg, col_reg}>=10'b1100000101) && ({row_reg, col_reg}<10'b1100001100)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}>=10'b1100001100) && ({row_reg, col_reg}<10'b1100001110)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}==10'b1100001110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100001111)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1100010000)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}>=10'b1100010001) && ({row_reg, col_reg}<10'b1100010011)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}>=10'b1100010011) && ({row_reg, col_reg}<10'b1100010110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100010110)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1100010111) && ({row_reg, col_reg}<10'b1100011011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100011011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b1100011100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b1100011101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1100100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b1100100001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1100100010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}>=10'b1100100011) && ({row_reg, col_reg}<10'b1100100101)) color_data = 12'b110100110110;
		if(({row_reg, col_reg}==10'b1100100101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100100110)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1100100111) && ({row_reg, col_reg}<10'b1100101111)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100101111)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1100110000) && ({row_reg, col_reg}<10'b1100110101)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100110101)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1100110110) && ({row_reg, col_reg}<10'b1100111011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1100111011)) color_data = 12'b110000010100;
		if(({row_reg, col_reg}==10'b1100111100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b1100111101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1101000000)) color_data = 12'b111010001010;
		if(({row_reg, col_reg}==10'b1101000001)) color_data = 12'b111110011011;
		if(({row_reg, col_reg}==10'b1101000010)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b1101000011)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}==10'b1101000100)) color_data = 12'b110101000110;
		if(({row_reg, col_reg}>=10'b1101000101) && ({row_reg, col_reg}<10'b1101001000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1101001000)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}==10'b1101001001)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1101001010)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1101001011) && ({row_reg, col_reg}<10'b1101010000)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1101010000)) color_data = 12'b111001000110;
		if(({row_reg, col_reg}>=10'b1101010001) && ({row_reg, col_reg}<10'b1101010011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1101010011)) color_data = 12'b111100110110;
		if(({row_reg, col_reg}>=10'b1101010100) && ({row_reg, col_reg}<10'b1101010110)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1101010110)) color_data = 12'b111001000111;
		if(({row_reg, col_reg}>=10'b1101010111) && ({row_reg, col_reg}<10'b1101011001)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}>=10'b1101011001) && ({row_reg, col_reg}<10'b1101011011)) color_data = 12'b111000110110;
		if(({row_reg, col_reg}==10'b1101011011)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==10'b1101011100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b1101011101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1101100000)) color_data = 12'b111110001010;
		if(({row_reg, col_reg}==10'b1101100001)) color_data = 12'b111101111001;
		if(({row_reg, col_reg}==10'b1101100010)) color_data = 12'b110001000111;
		if(({row_reg, col_reg}==10'b1101100011)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}>=10'b1101100100) && ({row_reg, col_reg}<10'b1101100110)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}>=10'b1101100110) && ({row_reg, col_reg}<10'b1101101100)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}>=10'b1101101100) && ({row_reg, col_reg}<10'b1101101111)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b1101101111)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==10'b1101110000)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b1101110001)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==10'b1101110010)) color_data = 12'b110100010101;
		if(({row_reg, col_reg}>=10'b1101110011) && ({row_reg, col_reg}<10'b1101110101)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}>=10'b1101110101) && ({row_reg, col_reg}<10'b1101111000)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b1101111000)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}>=10'b1101111001) && ({row_reg, col_reg}<10'b1101111011)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==10'b1101111011)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==10'b1101111100)) color_data = 12'b101000100100;

		if(({row_reg, col_reg}==10'b1101111101)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1110000000)) color_data = 12'b111001011000;
		if(({row_reg, col_reg}==10'b1110000001)) color_data = 12'b110101000111;
		if(({row_reg, col_reg}>=10'b1110000010) && ({row_reg, col_reg}<10'b1110000110)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1110000110)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}>=10'b1110000111) && ({row_reg, col_reg}<10'b1110010001)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1110010001)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==10'b1110010010)) color_data = 12'b110000010100;
		if(({row_reg, col_reg}==10'b1110010011)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}>=10'b1110010100) && ({row_reg, col_reg}<10'b1110011001)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}>=10'b1110011001) && ({row_reg, col_reg}<10'b1110011011)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}>=10'b1110011011) && ({row_reg, col_reg}<10'b1110011101)) color_data = 12'b100100010100;

		if(({row_reg, col_reg}==10'b1110011101)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==10'b1110100000)) color_data = 12'b110100100101;
		if(({row_reg, col_reg}==10'b1110100001)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==10'b1110100010)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==10'b1110100011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}>=10'b1110100100) && ({row_reg, col_reg}<10'b1110100110)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}>=10'b1110100110) && ({row_reg, col_reg}<10'b1110101111)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}>=10'b1110101111) && ({row_reg, col_reg}<10'b1110110001)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1110110001)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1110110010)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==10'b1110110011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}>=10'b1110110100) && ({row_reg, col_reg}<10'b1110111010)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==10'b1110111010)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==10'b1110111011)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==10'b1110111100)) color_data = 12'b100000010011;

		if(({row_reg, col_reg}>=10'b1110111101) && ({row_reg, col_reg}<=10'b1110111101)) color_data = 12'b011000000010;
	end
endmodule