module tile_rom_2
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}==10'b0000000000)) color_data = 12'b010001000010;
		if(({row_reg, col_reg}==10'b0000000001)) color_data = 12'b110011001010;
		if(({row_reg, col_reg}==10'b0000000010)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b0000000011)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0000000100)) color_data = 12'b111011111100;
		if(({row_reg, col_reg}==10'b0000000101)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==10'b0000000110)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}>=10'b0000000111) && ({row_reg, col_reg}<10'b0000001001)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b0000001001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}>=10'b0000001010) && ({row_reg, col_reg}<10'b0000001100)) color_data = 12'b111011111110;
		if(({row_reg, col_reg}==10'b0000001100)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=10'b0000001101) && ({row_reg, col_reg}<10'b0000001111)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0000001111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==10'b0000010000)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0000010001)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==10'b0000010010)) color_data = 12'b110111111101;
		if(({row_reg, col_reg}==10'b0000010011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=10'b0000010100) && ({row_reg, col_reg}<10'b0000010110)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}>=10'b0000010110) && ({row_reg, col_reg}<10'b0000011000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=10'b0000011000) && ({row_reg, col_reg}<10'b0000011011)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}>=10'b0000011011) && ({row_reg, col_reg}<10'b0000011101)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}==10'b0000011101)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==10'b0000100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0000100001)) color_data = 12'b111011011100;
		if(({row_reg, col_reg}==10'b0000100010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}>=10'b0000100011) && ({row_reg, col_reg}<10'b0000101000)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}>=10'b0000101000) && ({row_reg, col_reg}<10'b0000101101)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}>=10'b0000101101) && ({row_reg, col_reg}<10'b0000101111)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0000101111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=10'b0000110000) && ({row_reg, col_reg}<10'b0000111001)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}>=10'b0000111001) && ({row_reg, col_reg}<10'b0000111101)) color_data = 12'b111111111101;

		if(({row_reg, col_reg}==10'b0000111101)) color_data = 12'b111011101011;
		if(({row_reg, col_reg}==10'b0001000000)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==10'b0001000001)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b0001000010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b0001000011)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==10'b0001000100)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0001000101)) color_data = 12'b110111011010;
		if(({row_reg, col_reg}==10'b0001000110)) color_data = 12'b110111101010;
		if(({row_reg, col_reg}==10'b0001000111)) color_data = 12'b111011101011;
		if(({row_reg, col_reg}==10'b0001001000)) color_data = 12'b110111101011;
		if(({row_reg, col_reg}==10'b0001001001)) color_data = 12'b111011011011;
		if(({row_reg, col_reg}>=10'b0001001010) && ({row_reg, col_reg}<10'b0001001100)) color_data = 12'b111111011011;
		if(({row_reg, col_reg}==10'b0001001100)) color_data = 12'b111111001011;
		if(({row_reg, col_reg}==10'b0001001101)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0001001110)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0001001111)) color_data = 12'b110111101010;
		if(({row_reg, col_reg}==10'b0001010000)) color_data = 12'b111111001010;
		if(({row_reg, col_reg}==10'b0001010001)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0001010010) && ({row_reg, col_reg}<10'b0001011000)) color_data = 12'b111011011011;
		if(({row_reg, col_reg}>=10'b0001011000) && ({row_reg, col_reg}<10'b0001011010)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0001011010)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0001011011)) color_data = 12'b111011101011;
		if(({row_reg, col_reg}==10'b0001011100)) color_data = 12'b110111001001;

		if(({row_reg, col_reg}==10'b0001011101)) color_data = 12'b110110111000;
		if(({row_reg, col_reg}==10'b0001100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0001100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0001100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0001100011)) color_data = 12'b111011001010;
		if(({row_reg, col_reg}==10'b0001100100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0001100101) && ({row_reg, col_reg}<10'b0001100111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0001100111) && ({row_reg, col_reg}<10'b0001101010)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0001101010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0001101011) && ({row_reg, col_reg}<10'b0001101110)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0001101110) && ({row_reg, col_reg}<10'b0001110000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0001110000) && ({row_reg, col_reg}<10'b0001110100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0001110100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0001110101) && ({row_reg, col_reg}<10'b0001110111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0001110111) && ({row_reg, col_reg}<10'b0001111010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0001111010) && ({row_reg, col_reg}<10'b0001111100)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0001111100)) color_data = 12'b110010110111;

		if(({row_reg, col_reg}==10'b0001111101)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b0010000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0010000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0010000010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b0010000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0010000100)) color_data = 12'b111111101011;
		if(({row_reg, col_reg}==10'b0010000101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010000110)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0010000111) && ({row_reg, col_reg}<10'b0010001001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010001001)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0010001010) && ({row_reg, col_reg}<10'b0010001101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0010001101) && ({row_reg, col_reg}<10'b0010010000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0010010000) && ({row_reg, col_reg}<10'b0010010011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010010011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0010010100) && ({row_reg, col_reg}<10'b0010010110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010010110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0010010111) && ({row_reg, col_reg}<10'b0010011010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010011010)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b0010011011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010011100)) color_data = 12'b110010100110;

		if(({row_reg, col_reg}==10'b0010011101)) color_data = 12'b110010010101;
		if(({row_reg, col_reg}==10'b0010100000)) color_data = 12'b100010010110;
		if(({row_reg, col_reg}==10'b0010100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0010100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0010100011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0010100100)) color_data = 12'b111111101011;
		if(({row_reg, col_reg}==10'b0010100101)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0010100110)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0010100111) && ({row_reg, col_reg}<10'b0010101100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010101100)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0010101101)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b0010101110) && ({row_reg, col_reg}<10'b0010110000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0010110000)) color_data = 12'b111011111001;
		if(({row_reg, col_reg}==10'b0010110001)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b0010110010) && ({row_reg, col_reg}<10'b0010111000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0010111000) && ({row_reg, col_reg}<10'b0010111011)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0010111011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0010111100)) color_data = 12'b110010100110;

		if(({row_reg, col_reg}==10'b0010111101)) color_data = 12'b110010100101;
		if(({row_reg, col_reg}==10'b0011000000)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==10'b0011000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0011000010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b0011000011)) color_data = 12'b111011001010;
		if(({row_reg, col_reg}==10'b0011000100)) color_data = 12'b111111101011;
		if(({row_reg, col_reg}==10'b0011000101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0011000110) && ({row_reg, col_reg}<10'b0011001000)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0011001000) && ({row_reg, col_reg}<10'b0011001011)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0011001011) && ({row_reg, col_reg}<10'b0011001101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0011001101)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0011001110) && ({row_reg, col_reg}<10'b0011010011)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b0011010011) && ({row_reg, col_reg}<10'b0011010110)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0011010110) && ({row_reg, col_reg}<10'b0011011000)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b0011011000) && ({row_reg, col_reg}<10'b0011011100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0011011100)) color_data = 12'b110010110110;

		if(({row_reg, col_reg}==10'b0011011101)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b0011100000)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==10'b0011100001)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==10'b0011100010)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0011100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0011100100)) color_data = 12'b111111101011;
		if(({row_reg, col_reg}>=10'b0011100101) && ({row_reg, col_reg}<10'b0011100111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0011100111) && ({row_reg, col_reg}<10'b0011101111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0011101111) && ({row_reg, col_reg}<10'b0011110001)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0011110001) && ({row_reg, col_reg}<10'b0011111000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0011111000)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0011111001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0011111010)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0011111011)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b0011111100) && ({row_reg, col_reg}<10'b0100000000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b0100000000)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==10'b0100000001)) color_data = 12'b111111111110;
		if(({row_reg, col_reg}==10'b0100000010)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b0100000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0100000100)) color_data = 12'b111011101011;
		if(({row_reg, col_reg}==10'b0100000101)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0100000110) && ({row_reg, col_reg}<10'b0100001000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0100001000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0100001001) && ({row_reg, col_reg}<10'b0100001100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0100001100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0100001101)) color_data = 12'b111110111001;
		if(({row_reg, col_reg}>=10'b0100001110) && ({row_reg, col_reg}<10'b0100010001)) color_data = 12'b111110000110;
		if(({row_reg, col_reg}==10'b0100010001)) color_data = 12'b111110100111;
		if(({row_reg, col_reg}==10'b0100010010)) color_data = 12'b111111011001;
		if(({row_reg, col_reg}>=10'b0100010011) && ({row_reg, col_reg}<10'b0100011100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0100011100)) color_data = 12'b110010100111;

		if(({row_reg, col_reg}==10'b0100011101)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b0100100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==10'b0100100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0100100010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b0100100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0100100100)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0100100101) && ({row_reg, col_reg}<10'b0100101000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0100101000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0100101001) && ({row_reg, col_reg}<10'b0100101011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0100101011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0100101100)) color_data = 12'b111010010111;
		if(({row_reg, col_reg}==10'b0100101101)) color_data = 12'b110001010011;
		if(({row_reg, col_reg}==10'b0100101110)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b0100101111)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b0100110000)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b0100110001)) color_data = 12'b110001010011;
		if(({row_reg, col_reg}==10'b0100110010)) color_data = 12'b110101110101;
		if(({row_reg, col_reg}==10'b0100110011)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}>=10'b0100110100) && ({row_reg, col_reg}<10'b0100111100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0100111100)) color_data = 12'b110110100111;

		if(({row_reg, col_reg}==10'b0100111101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b0101000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0101000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0101000010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b0101000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b0101000100) && ({row_reg, col_reg}<10'b0101000110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0101000110) && ({row_reg, col_reg}<10'b0101001001)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0101001001) && ({row_reg, col_reg}<10'b0101001011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0101001011)) color_data = 12'b111110100111;
		if(({row_reg, col_reg}>=10'b0101001100) && ({row_reg, col_reg}<10'b0101001110)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b0101001110)) color_data = 12'b111001110110;
		if(({row_reg, col_reg}==10'b0101001111)) color_data = 12'b111010010110;
		if(({row_reg, col_reg}==10'b0101010000)) color_data = 12'b111010000110;
		if(({row_reg, col_reg}==10'b0101010001)) color_data = 12'b110101100100;
		if(({row_reg, col_reg}==10'b0101010010)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b0101010011)) color_data = 12'b111010000101;
		if(({row_reg, col_reg}==10'b0101010100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0101010101) && ({row_reg, col_reg}<10'b0101010111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0101010111)) color_data = 12'b111111011001;
		if(({row_reg, col_reg}>=10'b0101011000) && ({row_reg, col_reg}<10'b0101011010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0101011010)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0101011011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0101011100)) color_data = 12'b110110100110;

		if(({row_reg, col_reg}==10'b0101011101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b0101100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0101100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0101100010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b0101100011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b0101100100) && ({row_reg, col_reg}<10'b0101100110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0101100110) && ({row_reg, col_reg}<10'b0101101001)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0101101001)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b0101101010)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0101101011)) color_data = 12'b110110000101;
		if(({row_reg, col_reg}==10'b0101101100)) color_data = 12'b110001000011;
		if(({row_reg, col_reg}==10'b0101101101)) color_data = 12'b111110010111;
		if(({row_reg, col_reg}==10'b0101101110)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}>=10'b0101101111) && ({row_reg, col_reg}<10'b0101110001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0101110001)) color_data = 12'b111110100111;
		if(({row_reg, col_reg}==10'b0101110010)) color_data = 12'b111001010011;
		if(({row_reg, col_reg}==10'b0101110011)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b0101110100)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b0101110101)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0101110110)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0101110111)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0101111000) && ({row_reg, col_reg}<10'b0101111100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0101111100)) color_data = 12'b110010100110;

		if(({row_reg, col_reg}==10'b0101111101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b0110000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0110000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0110000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0110000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b0110000100) && ({row_reg, col_reg}<10'b0110000110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0110000110) && ({row_reg, col_reg}<10'b0110001000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0110001000)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0110001001)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b0110001010)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0110001011)) color_data = 12'b111010100111;
		if(({row_reg, col_reg}==10'b0110001100)) color_data = 12'b111010010110;
		if(({row_reg, col_reg}==10'b0110001101)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}>=10'b0110001110) && ({row_reg, col_reg}<10'b0110010000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0110010000)) color_data = 12'b110111111010;
		if(({row_reg, col_reg}==10'b0110010001)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b0110010010)) color_data = 12'b111101100100;
		if(({row_reg, col_reg}==10'b0110010011)) color_data = 12'b111001010011;
		if(({row_reg, col_reg}==10'b0110010100)) color_data = 12'b111110111000;
		if(({row_reg, col_reg}==10'b0110010101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0110010110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0110010111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0110011000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0110011001) && ({row_reg, col_reg}<10'b0110011100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b0110011100) && ({row_reg, col_reg}<10'b0110100000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b0110100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0110100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0110100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0110100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b0110100100) && ({row_reg, col_reg}<10'b0110101000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0110101000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0110101001) && ({row_reg, col_reg}<10'b0110110000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0110110000)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0110110001)) color_data = 12'b111110111000;
		if(({row_reg, col_reg}==10'b0110110010)) color_data = 12'b111001010100;
		if(({row_reg, col_reg}==10'b0110110011)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b0110110100)) color_data = 12'b111111001000;
		if(({row_reg, col_reg}==10'b0110110101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0110110110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0110110111)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0110111000) && ({row_reg, col_reg}<10'b0110111100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b0110111100) && ({row_reg, col_reg}<10'b0111000000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b0111000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b0111000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0111000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b0111000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0111000100)) color_data = 12'b111111101011;
		if(({row_reg, col_reg}>=10'b0111000101) && ({row_reg, col_reg}<10'b0111000111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0111000111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111001000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0111001001) && ({row_reg, col_reg}<10'b0111001101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111001101)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b0111001110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111001111)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0111010000)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b0111010001)) color_data = 12'b111001110101;
		if(({row_reg, col_reg}==10'b0111010010)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b0111010011)) color_data = 12'b110101100100;
		if(({row_reg, col_reg}==10'b0111010100)) color_data = 12'b111111011001;
		if(({row_reg, col_reg}==10'b0111010101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111010110)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0111010111)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b0111011000) && ({row_reg, col_reg}<10'b0111011100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111011100)) color_data = 12'b110010100110;

		if(({row_reg, col_reg}==10'b0111011101)) color_data = 12'b101110100110;
		if(({row_reg, col_reg}==10'b0111100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==10'b0111100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b0111100010)) color_data = 12'b111111101101;
		if(({row_reg, col_reg}==10'b0111100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b0111100100)) color_data = 12'b111011101011;
		if(({row_reg, col_reg}==10'b0111100101)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==10'b0111100110)) color_data = 12'b110111111010;
		if(({row_reg, col_reg}==10'b0111100111)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==10'b0111101000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b0111101001) && ({row_reg, col_reg}<10'b0111101100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b0111101100)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b0111101101)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b0111101110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111101111)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b0111110000)) color_data = 12'b111101110110;
		if(({row_reg, col_reg}==10'b0111110001)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b0111110010)) color_data = 12'b110101010100;
		if(({row_reg, col_reg}==10'b0111110011)) color_data = 12'b111110101000;
		if(({row_reg, col_reg}==10'b0111110100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111110101)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b0111110110) && ({row_reg, col_reg}<10'b0111111100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b0111111100)) color_data = 12'b110010100111;

		if(({row_reg, col_reg}==10'b0111111101)) color_data = 12'b101110100110;
		if(({row_reg, col_reg}==10'b1000000000)) color_data = 12'b011110010110;
		if(({row_reg, col_reg}==10'b1000000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1000000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1000000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b1000000100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b1000000101) && ({row_reg, col_reg}<10'b1000001101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1000001101) && ({row_reg, col_reg}<10'b1000001111)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1000001111)) color_data = 12'b111010000101;
		if(({row_reg, col_reg}==10'b1000010000)) color_data = 12'b111001010011;
		if(({row_reg, col_reg}==10'b1000010001)) color_data = 12'b110001010011;
		if(({row_reg, col_reg}==10'b1000010010)) color_data = 12'b111110100111;
		if(({row_reg, col_reg}==10'b1000010011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000010100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b1000010101) && ({row_reg, col_reg}<10'b1000010111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000010111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1000011000)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==10'b1000011001)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1000011010) && ({row_reg, col_reg}<10'b1000011100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000011100)) color_data = 12'b110110100110;

		if(({row_reg, col_reg}==10'b1000011101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b1000100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1000100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1000100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1000100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b1000100100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b1000100101) && ({row_reg, col_reg}<10'b1000100111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000100111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1000101000)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b1000101001) && ({row_reg, col_reg}<10'b1000101101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000101101)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1000101110)) color_data = 12'b110110000110;
		if(({row_reg, col_reg}==10'b1000101111)) color_data = 12'b110001100011;
		if(({row_reg, col_reg}==10'b1000110000)) color_data = 12'b101101100011;
		if(({row_reg, col_reg}==10'b1000110001)) color_data = 12'b111010111000;
		if(({row_reg, col_reg}>=10'b1000110010) && ({row_reg, col_reg}<10'b1000110110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000110110)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b1000110111) && ({row_reg, col_reg}<10'b1000111001)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1000111001) && ({row_reg, col_reg}<10'b1000111100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1000111100)) color_data = 12'b110110100110;

		if(({row_reg, col_reg}==10'b1000111101)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b1001000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1001000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1001000010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b1001000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1001000100) && ({row_reg, col_reg}<10'b1001000111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001000111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1001001000)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b1001001001)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==10'b1001001010)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1001001011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001001100)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1001001101)) color_data = 12'b110110000110;
		if(({row_reg, col_reg}==10'b1001001110)) color_data = 12'b101101010011;
		if(({row_reg, col_reg}==10'b1001001111)) color_data = 12'b110101100100;
		if(({row_reg, col_reg}==10'b1001010000)) color_data = 12'b110110111000;
		if(({row_reg, col_reg}>=10'b1001010001) && ({row_reg, col_reg}<10'b1001010011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1001010011) && ({row_reg, col_reg}<10'b1001010101)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1001010101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001010110)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}>=10'b1001010111) && ({row_reg, col_reg}<10'b1001011100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b1001011100) && ({row_reg, col_reg}<10'b1001100000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b1001100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1001100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1001100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1001100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1001100100) && ({row_reg, col_reg}<10'b1001101000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001101000)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b1001101001) && ({row_reg, col_reg}<10'b1001101011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001101011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1001101100)) color_data = 12'b111010000110;
		if(({row_reg, col_reg}==10'b1001101101)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b1001101110)) color_data = 12'b111001010011;
		if(({row_reg, col_reg}==10'b1001101111)) color_data = 12'b111110000111;
		if(({row_reg, col_reg}>=10'b1001110000) && ({row_reg, col_reg}<10'b1001110011)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b1001110011)) color_data = 12'b111111011001;
		if(({row_reg, col_reg}==10'b1001110100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001110101)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b1001110110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1001110111)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b1001111000) && ({row_reg, col_reg}<10'b1001111100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b1001111100) && ({row_reg, col_reg}<10'b1010000000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b1010000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1010000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1010000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1010000011)) color_data = 12'b110111011010;
		if(({row_reg, col_reg}>=10'b1010000100) && ({row_reg, col_reg}<10'b1010000110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1010000110) && ({row_reg, col_reg}<10'b1010001010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1010001010)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1010001011)) color_data = 12'b111010000110;
		if(({row_reg, col_reg}==10'b1010001100)) color_data = 12'b110101000011;
		if(({row_reg, col_reg}==10'b1010001101)) color_data = 12'b111101000100;
		if(({row_reg, col_reg}>=10'b1010001110) && ({row_reg, col_reg}<10'b1010010000)) color_data = 12'b111101000011;
		if(({row_reg, col_reg}>=10'b1010010000) && ({row_reg, col_reg}<10'b1010010010)) color_data = 12'b111001010100;
		if(({row_reg, col_reg}==10'b1010010010)) color_data = 12'b111001100100;
		if(({row_reg, col_reg}==10'b1010010011)) color_data = 12'b110101110100;
		if(({row_reg, col_reg}==10'b1010010100)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b1010010101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1010010110)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b1010010111) && ({row_reg, col_reg}<10'b1010011100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b1010011100) && ({row_reg, col_reg}<10'b1010100000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b1010100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1010100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1010100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1010100011)) color_data = 12'b110111011010;
		if(({row_reg, col_reg}>=10'b1010100100) && ({row_reg, col_reg}<10'b1010100110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1010100110) && ({row_reg, col_reg}<10'b1010101000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1010101000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b1010101001) && ({row_reg, col_reg}<10'b1010101011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1010101011)) color_data = 12'b110110000101;
		if(({row_reg, col_reg}==10'b1010101100)) color_data = 12'b110101100100;
		if(({row_reg, col_reg}==10'b1010101101)) color_data = 12'b111001010011;
		if(({row_reg, col_reg}==10'b1010101110)) color_data = 12'b111001010100;
		if(({row_reg, col_reg}>=10'b1010101111) && ({row_reg, col_reg}<10'b1010110010)) color_data = 12'b110101010011;
		if(({row_reg, col_reg}==10'b1010110010)) color_data = 12'b111001010100;
		if(({row_reg, col_reg}==10'b1010110011)) color_data = 12'b110001100011;
		if(({row_reg, col_reg}==10'b1010110100)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}>=10'b1010110101) && ({row_reg, col_reg}<10'b1010111100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b1010111100) && ({row_reg, col_reg}<10'b1011000000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b1011000000)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==10'b1011000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1011000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1011000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1011000100) && ({row_reg, col_reg}<10'b1011000110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1011000110) && ({row_reg, col_reg}<10'b1011001001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011001001)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b1011001010)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b1011001011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}>=10'b1011001100) && ({row_reg, col_reg}<10'b1011001111)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b1011001111)) color_data = 12'b111111011001;
		if(({row_reg, col_reg}>=10'b1011010000) && ({row_reg, col_reg}<10'b1011010100)) color_data = 12'b111111001001;
		if(({row_reg, col_reg}==10'b1011010100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1011010101) && ({row_reg, col_reg}<10'b1011011000)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}>=10'b1011011000) && ({row_reg, col_reg}<10'b1011011100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011011100)) color_data = 12'b110010100110;

		if(({row_reg, col_reg}==10'b1011011101)) color_data = 12'b101110100110;
		if(({row_reg, col_reg}==10'b1011100000)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==10'b1011100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1011100010)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b1011100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1011100100) && ({row_reg, col_reg}<10'b1011101001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011101001)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b1011101010)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}>=10'b1011101011) && ({row_reg, col_reg}<10'b1011101101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011101101)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b1011101110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011101111)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1011110000)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==10'b1011110001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011110010)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1011110011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1011110100)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1011110101)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b1011110110) && ({row_reg, col_reg}<10'b1011111100)) color_data = 12'b111111101010;

		if(({row_reg, col_reg}>=10'b1011111100) && ({row_reg, col_reg}<10'b1100000000)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}==10'b1100000000)) color_data = 12'b100110000110;
		if(({row_reg, col_reg}==10'b1100000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1100000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1100000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1100000100) && ({row_reg, col_reg}<10'b1100001100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1100001100) && ({row_reg, col_reg}<10'b1100010000)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1100010000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1100010001) && ({row_reg, col_reg}<10'b1100011001)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1100011001) && ({row_reg, col_reg}<10'b1100011100)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1100011100)) color_data = 12'b110110100111;

		if(({row_reg, col_reg}==10'b1100011101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b1100100000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1100100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1100100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1100100011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1100100100) && ({row_reg, col_reg}<10'b1100100110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1100100110)) color_data = 12'b111111101001;
		if(({row_reg, col_reg}==10'b1100100111)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}>=10'b1100101000) && ({row_reg, col_reg}<10'b1100101101)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1100101101)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1100101110) && ({row_reg, col_reg}<10'b1100110011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1100110011)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1100110100) && ({row_reg, col_reg}<10'b1100110111)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1100110111)) color_data = 12'b111011111010;
		if(({row_reg, col_reg}==10'b1100111000)) color_data = 12'b111011101001;
		if(({row_reg, col_reg}==10'b1100111001)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b1100111010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1100111011)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1100111100)) color_data = 12'b110110100110;

		if(({row_reg, col_reg}==10'b1100111101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b1101000000)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==10'b1101000001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1101000010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1101000011)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}>=10'b1101000100) && ({row_reg, col_reg}<10'b1101000110)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1101000110) && ({row_reg, col_reg}<10'b1101001000)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}>=10'b1101001000) && ({row_reg, col_reg}<10'b1101001010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1101001010)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1101001011)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1101001100) && ({row_reg, col_reg}<10'b1101001110)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1101001110) && ({row_reg, col_reg}<10'b1101010000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1101010000)) color_data = 12'b111111011010;
		if(({row_reg, col_reg}==10'b1101010001)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}>=10'b1101010010) && ({row_reg, col_reg}<10'b1101010100)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}>=10'b1101010100) && ({row_reg, col_reg}<10'b1101011000)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1101011000)) color_data = 12'b111011101010;
		if(({row_reg, col_reg}==10'b1101011001)) color_data = 12'b111111111010;
		if(({row_reg, col_reg}==10'b1101011010)) color_data = 12'b111111101010;
		if(({row_reg, col_reg}==10'b1101011011)) color_data = 12'b111111011001;

		if(({row_reg, col_reg}>=10'b1101011100) && ({row_reg, col_reg}<10'b1101100000)) color_data = 12'b110110100110;
		if(({row_reg, col_reg}==10'b1101100000)) color_data = 12'b100010010110;
		if(({row_reg, col_reg}==10'b1101100001)) color_data = 12'b111111111101;
		if(({row_reg, col_reg}==10'b1101100010)) color_data = 12'b111111111100;
		if(({row_reg, col_reg}==10'b1101100011)) color_data = 12'b110111001001;
		if(({row_reg, col_reg}>=10'b1101100100) && ({row_reg, col_reg}<10'b1101100110)) color_data = 12'b110111001000;
		if(({row_reg, col_reg}==10'b1101100110)) color_data = 12'b110111000111;
		if(({row_reg, col_reg}>=10'b1101100111) && ({row_reg, col_reg}<10'b1101101001)) color_data = 12'b110111001000;
		if(({row_reg, col_reg}>=10'b1101101001) && ({row_reg, col_reg}<10'b1101101011)) color_data = 12'b111011001000;
		if(({row_reg, col_reg}>=10'b1101101011) && ({row_reg, col_reg}<10'b1101101111)) color_data = 12'b110111001000;
		if(({row_reg, col_reg}>=10'b1101101111) && ({row_reg, col_reg}<10'b1101110001)) color_data = 12'b111011001000;
		if(({row_reg, col_reg}>=10'b1101110001) && ({row_reg, col_reg}<10'b1101110100)) color_data = 12'b110111001000;
		if(({row_reg, col_reg}==10'b1101110100)) color_data = 12'b111011001000;
		if(({row_reg, col_reg}==10'b1101110101)) color_data = 12'b111010111000;
		if(({row_reg, col_reg}>=10'b1101110110) && ({row_reg, col_reg}<10'b1101111000)) color_data = 12'b111011001000;
		if(({row_reg, col_reg}==10'b1101111000)) color_data = 12'b110111000111;
		if(({row_reg, col_reg}==10'b1101111001)) color_data = 12'b111011001000;
		if(({row_reg, col_reg}>=10'b1101111010) && ({row_reg, col_reg}<10'b1101111100)) color_data = 12'b111010111000;
		if(({row_reg, col_reg}==10'b1101111100)) color_data = 12'b110010010110;

		if(({row_reg, col_reg}==10'b1101111101)) color_data = 12'b110010010101;
		if(({row_reg, col_reg}==10'b1110000000)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==10'b1110000001)) color_data = 12'b111111101100;
		if(({row_reg, col_reg}==10'b1110000010)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b1110000011)) color_data = 12'b110010110111;
		if(({row_reg, col_reg}==10'b1110000100)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}>=10'b1110000101) && ({row_reg, col_reg}<10'b1110000111)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==10'b1110000111)) color_data = 12'b101110100101;
		if(({row_reg, col_reg}==10'b1110001000)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==10'b1110001001)) color_data = 12'b110010010101;
		if(({row_reg, col_reg}==10'b1110001010)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}>=10'b1110001011) && ({row_reg, col_reg}<10'b1110001110)) color_data = 12'b101110010110;
		if(({row_reg, col_reg}==10'b1110001110)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b1110001111)) color_data = 12'b110010010101;
		if(({row_reg, col_reg}>=10'b1110010000) && ({row_reg, col_reg}<10'b1110010010)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b1110010010)) color_data = 12'b101110010110;
		if(({row_reg, col_reg}==10'b1110010011)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}>=10'b1110010100) && ({row_reg, col_reg}<10'b1110011011)) color_data = 12'b110010010101;
		if(({row_reg, col_reg}==10'b1110011011)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==10'b1110011100)) color_data = 12'b101110010101;

		if(({row_reg, col_reg}==10'b1110011101)) color_data = 12'b101010000100;
		if(({row_reg, col_reg}==10'b1110100000)) color_data = 12'b011101110100;
		if(({row_reg, col_reg}==10'b1110100001)) color_data = 12'b111011011010;
		if(({row_reg, col_reg}==10'b1110100010)) color_data = 12'b110111001001;
		if(({row_reg, col_reg}>=10'b1110100011) && ({row_reg, col_reg}<10'b1110100101)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}>=10'b1110100101) && ({row_reg, col_reg}<10'b1110101001)) color_data = 12'b110110100110;
		if(({row_reg, col_reg}>=10'b1110101001) && ({row_reg, col_reg}<10'b1110101011)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}>=10'b1110101011) && ({row_reg, col_reg}<10'b1110101101)) color_data = 12'b110110100110;
		if(({row_reg, col_reg}>=10'b1110101101) && ({row_reg, col_reg}<10'b1110110101)) color_data = 12'b110110010110;
		if(({row_reg, col_reg}>=10'b1110110101) && ({row_reg, col_reg}<10'b1110111001)) color_data = 12'b110110100110;
		if(({row_reg, col_reg}==10'b1110111001)) color_data = 12'b110010100110;
		if(({row_reg, col_reg}>=10'b1110111010) && ({row_reg, col_reg}<10'b1110111100)) color_data = 12'b110110100110;
		if(({row_reg, col_reg}==10'b1110111100)) color_data = 12'b110010100110;

		if(({row_reg, col_reg}>=10'b1110111101) && ({row_reg, col_reg}<=10'b1110111101)) color_data = 12'b101110000100;
	end
endmodule